module ram_output;

	reg signed [18:0] mem [63:0];

endmodule